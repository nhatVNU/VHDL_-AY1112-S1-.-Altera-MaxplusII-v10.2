LIBRARY IEEE;
USE IEEE. STD_LOGIC_1164.ALL;
USE IEEE. STD_LOGIC_ARITH.ALL;
USE IEEE. STD_LOGIC_UNSIGNED.ALL;

ENTITY IC74LS283 IS

PORT(
	a: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	b: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	c0: IN STD_LOGIC;
	s: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	c4: out STD_LOGIC
	);
END IC74LS283;

ARCHITECTURE behavior OF IC74LS283 IS

	SIGNAL a_temp: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL b_temp: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL sum_temp: STD_LOGIC_VECTOR (4 DOWNTO 0);
BEGIN
	a_temp <= '0'&a;
	b_temp <= '0'&b;
	sum_temp <= a_temp + b_temp+c0;
	
	s <= sum_temp(3 DOWNTO 0);
	c4 <= sum_temp(4);
END behavior;




LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY tn10 IS
PORT (
a, b : IN STD_LOGIC_VECTOR(3 downto 0);
d : OUT STD_LOGIC_VECTOR(3 downto 0);
c4: OUT STD_LOGIC);
END tn10;


ARCHITECTURE Structure OF tn10 IS
SIGNAL c : STD_LOGIC_VECTOR(1 to 3);
SIGNAL f : STD_LOGIC_VECTOR(3 downto 0);
SIGNAL c0: STD_LOGIC;
COMPONENT IC74LS283
PORT(
	a: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	b: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	c0: IN STD_LOGIC;
	s: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	c4: out STD_LOGIC
	);
END COMPONENT;

BEGIN
c0 <= '1';
f <= not b;
u0: IC74LS283 PORT MAP(a,f,c0,d,c4) ;

END Structure;
