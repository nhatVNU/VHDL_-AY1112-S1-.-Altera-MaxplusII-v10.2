LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY D_FF IS
PORT(
	D, CLK, PR, CL: IN STD_LOGIC;
	Q, Qn: BUFFER STD_LOGIC
);
END D_FF;
ARCHITECTURE BEHAVIOR OF D_FF IS
BEGIN 
	PROCESS(CLK, PR, CL)
	BEGIN	
		IF PR='0' THEN Q <= '1'; Qn <='0';
		ELSIF CL='0' THEN Q <= '0'; Qn <='1';
		ELSIF falling_edge(CLK) THEN Q <= D; Qn <= NOT Q;
	END IF;
	END PROCESS;
END BEHAVIOR;