LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY tn7 IS
	PORT ( c, b, a : IN STD_LOGIC;
	e,e1,e2: IN STD_LOGIC;
	y : OUT STD_LOGIC_VECTOR(7 downto 0));
END tn7;

ARCHITECTURE flow OF tn7 IS
SIGNAL data: STD_LOGIC_VECTOR(2 downto 0);
SIGNAL temp: STD_LOGIC_VECTOR(7 downto 0);
BEGIN
data <= c & b & a;
WITH data SELECT temp <= "11111110" WHEN "000" ,
"11111101" WHEN "001" ,
"11111011" WHEN "010" ,
"11110111" WHEN "011" ,
"11101111" WHEN "100" ,
"11011111" WHEN "101" ,
"10111111" WHEN "110" ,
"01111111" WHEN "111" ;
y <= temp WHEN (e AND NOT e1 AND NOT e2) = '1' 
ELSE "11111111"; 
END flow;